-- vga_adapter.vhd
-- Created on: Sa 9. Dez 09:07:21 CET 2023
-- Author(s): Yannick Reiß
-- Content:  Entity vga_adapter
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

